// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: upstream_monitor.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Thu Feb 18 07:48:09 2021
//=============================================================================
// Description: Monitor for upstream
//=============================================================================

`ifndef UPSTREAM_MONITOR_SV
`define UPSTREAM_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file upstream.tpl

class upstream_monitor extends uvm_monitor;

  `uvm_component_utils(upstream_monitor)

  virtual upstream_if vif;

  upstream_config     m_config;

  uvm_analysis_port #(ustream_trans) analysis_port;

  ustream_trans m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file upstream.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file upstream.tpl

endclass : upstream_monitor 


function upstream_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task upstream_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = ustream_trans::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file generated_tb/tb/include/upstream_monitor_inc.sv
task upstream_monitor::do_mon;
  forever @(vif.ustream_if.clk)
  begin
    m_trans.rand_instruction <= vif.ustream_if.lane0_txdata;
    `uvm_info(get_type_name(), $sformatf("txdata0: %X", vif.ustream_if.lane0_txdata), UVM_MEDIUM);
  end
endtask

// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file upstream.tpl

`endif // UPSTREAM_MONITOR_SV

