package verif_pkg;

  import dw_vip_pcie_uvm_pkg::*;

endpackage

