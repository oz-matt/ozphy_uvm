// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: downstream_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Wed Feb 17 10:05:16 2021
//=============================================================================
// Description: Sequencer for downstream
//=============================================================================

`ifndef DOWNSTREAM_SEQUENCER_SV
`define DOWNSTREAM_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(ustream_trans) downstream_sequencer_t;


`endif // DOWNSTREAM_SEQUENCER_SV

